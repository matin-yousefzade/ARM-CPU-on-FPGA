module Instruction_Memory (rst, address, readData);
  
  input [31:0] address;
  input rst;
  output [31:0] readData;
  
  reg [31:0] array [0:255];
  wire [7:0] index = address[31:2];
  integer i;
  
  assign readData = array[index];
   
  always @(posedge rst) begin
    for(i = 0; i < 256; i = i + 1) array[i] <= 32'h0;
    /*array[0] <= {4'b1110, 2'b00, 1'b1, 4'b1111, 1'b0, 4'h0, 4'h1, 12'hAB};
    array[1] <= {4'b1110, 2'b00, 1'b1, 4'b1101, 1'b0, 4'h0, 4'h2, 12'hAB};
    array[2] <= {4'b1110, 2'b01, 1'b0, 4'b0100, 1'b0, 4'h0, 4'h1, 12'h400};
    array[3] <= {4'b1110, 2'b01, 1'b0, 4'b0100, 1'b0, 4'h0, 4'h2, 12'h404};
    array[4] <= {4'b1110, 2'b01, 1'b0, 4'b0100, 1'b1, 4'h0, 4'h3, 12'h400};*/
    array[0] <= {32'b11100011101000000000000000010100}; //MOV R0 ,#20 //R0 = 20
    array[1] <= {32'b11100011101000000001101000000001}; //MOV R1 ,#4096 //R1 = 4096
    array[2] <= {32'b11100011101000000010000100000011}; //MOV R2 ,#0xC0000000 //R2 = -1073741824
    array[3] <= {32'b11100000100100100011000000000010}; //ADDS R3 ,R2,R2 //R3 = -2147483648
  	 array[4] <= {32'b11100000101000000100000000000000}; //ADC R4 ,R0,R0 //R4 = 41
    array[5] <= {32'b11100000010001000101000100000100}; //SUB R5 ,R4,R4,LSL #2 //R5 = -123
    array[6] <= {32'b11100000110000000110000010100000}; //SBC R6 ,R0,R0,LSR #1 //R6 = 9
    array[7] <= {32'b11100001100001010111000101000010}; //ORR R7 ,R5,R2,ASR #2 //R7 = -123
    array[8] <= {32'b11100000000001111000000000000011}; //AND R8 ,R7,R3 //R8 = -2147483648
    array[9] <= {32'b11100001111000001001000000000110}; //MVN R9 ,R6 //R9 = 10
    array[10] <= {32'b11100000001001001010000000000101}; //EOR R10,R4,R5 //R10 = -84
    array[11] <= {32'b11100001010110000000000000000110}; //CMP R8 ,R6
    array[12] <= {32'b00010000100000010001000000000001}; //ADDNE R1 ,R1,R1 //R1 = 8192
    array[13] <= {32'b11100001000110010000000000001000}; //TST R9 ,R8
    array[14] <= {32'b00000000100000100010000000000010}; //ADDEQ R2 ,R2,R2 //R2 = -1073741824
    array[15] <= {32'b11100011101000000000101100000001}; //MOV R0 ,#1024 //R0 = 1024
    array[16] <= {32'b11100100100000000001000000000000}; //STR R1 ,[R0],#0 //MEM[1024] = 8192
    array[17] <= {32'b11100100100100001011000000000000}; //LDR R11,[R0],#0 //R11 = 8192
    array[18] <= {32'b11100100100000000010000000000100}; //STR R2 ,[R0],#4 //MEM[1028] = -1073741824
    array[19] <= {32'b11100100100000000011000000001000}; //STR R3 ,[R0],#8 //MEM[1032] = -2147483648
    array[20] <= {32'b11100100100000000100000000001101}; //STR R4 ,[R0],#13 //MEM[1036] = 41
    array[21] <= {32'b11100100100000000101000000010000}; //STR R5 ,[R0],#16 //MEM[1040] = -123
    array[22] <= {32'b11100100100000000110000000010100}; //STR R6 ,[R0],#20 //MEM[1044] = 9
    array[23] <= {32'b11100100100100001010000000000100}; //LDR R10,[R0],#4 //R10 = -1073741824
    array[24] <= {32'b11100100100000000111000000011000}; //STR R7 ,[R0],#24 //MEM[1048] = -123
    array[25] <= {32'b11100011101000000001000000000100}; //MOV R1 ,#4 //R1 = 4
    array[26] <= {32'b11100011101000000010000000000000}; //MOV R2 ,#0 //R2 = 0
    array[27] <= {32'b11100011101000000011000000000000}; //MOV R3 ,#0 //R3 = 0
    array[28] <= {32'b11100000100000000100000100000011}; //ADD R4 ,R0,R3,LSL #2
    array[29] <= {32'b11100100100101000101000000000000}; //LDR R5 ,[R4],#0
    array[30] <= {32'b11100100100101000110000000000100}; //LDR R6 ,[R4],#4
    array[31] <= {32'b11100001010101010000000000000110}; //CMP R5 ,R6
    array[32] <= {32'b11000100100001000110000000000000}; //STRGT R6 ,[R4],#0
    array[33] <= {32'b11000100100001000101000000000100}; //STRGT R5 ,[R4],#4
    array[34] <= {32'b11100010100000110011000000000001}; //ADD R3 ,R3,#1
    array[35] <= {32'b11100011010100110000000000000011}; //CMP R3 ,#3
    array[36] <= {32'b10111010111111111111111111110111}; //BLT #-9
    array[37] <= {32'b11100010100000100010000000000001}; //ADD R2 ,R2,#1
    array[38] <= {32'b11100001010100100000000000000001}; //CMP R2 ,R1
    array[39] <= {32'b10111010111111111111111111110011}; //BLT #-13
    array[40] <= {32'b11100100100100000001000000000000}; //LDR R1 ,[R0],#0 //R1 = -2147483648
    array[41] <= {32'b11100100100100000010000000000100}; //LDR R2 ,[R0],#4 //R2 = -1073741824
    array[42] <= {32'b11100100100100000011000000001000}; //STR R3 ,[R0],#8 //R3 = 41
    array[43] <= {32'b11100100100100000100000000001100}; //STR R4 ,[R0],#12 //R4 = 8192
    array[44] <= {32'b11100100100100000101000000010000}; //STR R5 ,[R0],#16
    array[45] <= {32'b11100100100100000110000000010100}; //STR R6 ,[R0],#20
    array[46] <= {32'b11101010111111111111111111111111}; //B #-1
  end
  
endmodule